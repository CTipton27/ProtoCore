`timescale 1ns / 1ps
//FILE: sev_seg.v

module sev_seg(
    input clk,
    output [6:0] seg,
    output [1:0] an
    );
    
    wire[15:0] a;
    
endmodule
